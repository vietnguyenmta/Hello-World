use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
